library verilog;
use verilog.vl_types.all;
entity first_counter_tb is
end first_counter_tb;
